`timescale 1ns/1ns

module UART_Tx {
    parameter UART_CLK_CNT = 104;
}
{

}

endmodule